library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.VComponents.all;

entity patternMatch is
end patternMatch;

architecture Behavioral of patternMatch is

begin


end Behavioral;

